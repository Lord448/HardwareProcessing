-- NIOS2.vhd

-- Generated using ACDS version 22.1 922

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity NIOS2 is
	port (
		clk_clk                                       : in  std_logic                     := '0';             --                                    clk.clk
		control_pio_external_connection_export        : in  std_logic_vector(3 downto 0)  := (others => '0'); --        control_pio_external_connection.export
		dip_tx_data_pio_external_connection_export    : in  std_logic_vector(7 downto 0)  := (others => '0'); --    dip_tx_data_pio_external_connection.export
		parsedloop_irq_external_connection_export     : in  std_logic                     := '0';             --     parsedloop_irq_external_connection.export
		reset_reset_n                                 : in  std_logic                     := '0';             --                                  reset.reset_n
		start_timer_external_connection_export        : out std_logic;                                        --        start_timer_external_connection.export
		status_leds_pio_external_connection_export    : out std_logic_vector(3 downto 0);                     --    status_leds_pio_external_connection.export
		uart_rx_data_reg_external_connection_export   : in  std_logic_vector(7 downto 0)  := (others => '0'); --   uart_rx_data_reg_external_connection.export
		uart_rx_external_connection_export            : in  std_logic                     := '0';             --            uart_rx_external_connection.export
		uart_rx_pi_external_connection_export         : out std_logic_vector(31 downto 0);                    --         uart_rx_pi_external_connection.export
		uart_rx_status_reg_external_connection_export : in  std_logic_vector(1 downto 0)  := (others => '0'); -- uart_rx_status_reg_external_connection.export
		uart_tx_data_reg_external_connection_export   : out std_logic_vector(7 downto 0);                     --   uart_tx_data_reg_external_connection.export
		uart_tx_external_connection_export            : in  std_logic                     := '0';             --            uart_tx_external_connection.export
		uart_tx_po_external_connection_export         : out std_logic_vector(31 downto 0);                    --         uart_tx_po_external_connection.export
		uart_tx_start_external_connection_export      : out std_logic                                         --      uart_tx_start_external_connection.export
	);
end entity NIOS2;

architecture rtl of NIOS2 is
	component NIOS2_Control_PIO is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component NIOS2_Control_PIO;

	component NIOS2_DIP_TX_Data_PIO is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component NIOS2_DIP_TX_Data_PIO;

	component NIOS2_ParsedLoop_IRQ is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component NIOS2_ParsedLoop_IRQ;

	component NIOS2_Start_Timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component NIOS2_Start_Timer;

	component NIOS2_Status_LEDS_PIO is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component NIOS2_Status_LEDS_PIO;

	component NIOS2_UART_RX is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component NIOS2_UART_RX;

	component NIOS2_UART_RX_32_PO is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component NIOS2_UART_RX_32_PO;

	component NIOS2_UART_RX_STATUS_REG is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component NIOS2_UART_RX_STATUS_REG;

	component NIOS2_UART_TX_DATA_REG is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component NIOS2_UART_TX_DATA_REG;

	component NIOS2_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component NIOS2_jtag_uart_0;

	component NIOS2_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(15 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(15 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component NIOS2_nios2_gen2_0;

	component NIOS2_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component NIOS2_onchip_memory2_0;

	component NIOS2_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                  : in  std_logic                     := 'X';             -- clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_readdatavalid         : out std_logic;                                        -- readdatavalid
			nios2_gen2_0_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_instruction_master_readdatavalid  : out std_logic;                                        -- readdatavalid
			Control_PIO_s1_address                         : out std_logic_vector(2 downto 0);                     -- address
			Control_PIO_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DIP_TX_Data_PIO_s1_address                     : out std_logic_vector(1 downto 0);                     -- address
			DIP_TX_Data_PIO_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_address          : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write            : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read             : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write             : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read              : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                    : out std_logic_vector(11 downto 0);                    -- address
			onchip_memory2_0_s1_write                      : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                 : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                      : out std_logic;                                        -- clken
			ParsedLoop_IRQ_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			ParsedLoop_IRQ_s1_write                        : out std_logic;                                        -- write
			ParsedLoop_IRQ_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ParsedLoop_IRQ_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			ParsedLoop_IRQ_s1_chipselect                   : out std_logic;                                        -- chipselect
			Start_Timer_s1_address                         : out std_logic_vector(2 downto 0);                     -- address
			Start_Timer_s1_write                           : out std_logic;                                        -- write
			Start_Timer_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Start_Timer_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			Start_Timer_s1_chipselect                      : out std_logic;                                        -- chipselect
			Status_LEDS_PIO_s1_address                     : out std_logic_vector(2 downto 0);                     -- address
			Status_LEDS_PIO_s1_write                       : out std_logic;                                        -- write
			Status_LEDS_PIO_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Status_LEDS_PIO_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			Status_LEDS_PIO_s1_chipselect                  : out std_logic;                                        -- chipselect
			UART_RX_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			UART_RX_s1_write                               : out std_logic;                                        -- write
			UART_RX_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			UART_RX_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			UART_RX_s1_chipselect                          : out std_logic;                                        -- chipselect
			UART_RX_32_PO_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			UART_RX_32_PO_s1_write                         : out std_logic;                                        -- write
			UART_RX_32_PO_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			UART_RX_32_PO_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			UART_RX_32_PO_s1_chipselect                    : out std_logic;                                        -- chipselect
			UART_RX_DATA_REG_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			UART_RX_DATA_REG_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			UART_RX_STATUS_REG_s1_address                  : out std_logic_vector(1 downto 0);                     -- address
			UART_RX_STATUS_REG_s1_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			UART_TX_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			UART_TX_s1_write                               : out std_logic;                                        -- write
			UART_TX_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			UART_TX_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			UART_TX_s1_chipselect                          : out std_logic;                                        -- chipselect
			UART_TX_32_PO_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			UART_TX_32_PO_s1_write                         : out std_logic;                                        -- write
			UART_TX_32_PO_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			UART_TX_32_PO_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			UART_TX_32_PO_s1_chipselect                    : out std_logic;                                        -- chipselect
			UART_TX_DATA_REG_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			UART_TX_DATA_REG_s1_write                      : out std_logic;                                        -- write
			UART_TX_DATA_REG_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			UART_TX_DATA_REG_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			UART_TX_DATA_REG_s1_chipselect                 : out std_logic;                                        -- chipselect
			UART_TX_START_s1_address                       : out std_logic_vector(2 downto 0);                     -- address
			UART_TX_START_s1_write                         : out std_logic;                                        -- write
			UART_TX_START_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			UART_TX_START_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			UART_TX_START_s1_chipselect                    : out std_logic                                         -- chipselect
		);
	end component NIOS2_mm_interconnect_0;

	component NIOS2_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component NIOS2_irq_mapper;

	component nios2_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios2_rst_controller;

	component nios2_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component nios2_rst_controller_001;

	signal nios2_gen2_0_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                            : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                : std_logic_vector(15 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                   : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	signal nios2_gen2_0_data_master_write                                  : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                              : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                         : std_logic_vector(15 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                            : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal nios2_gen2_0_instruction_master_readdatavalid                   : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest      : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                  : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                   : std_logic_vector(11 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_uart_tx_32_po_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:UART_TX_32_PO_s1_chipselect -> UART_TX_32_PO:chipselect
	signal mm_interconnect_0_uart_tx_32_po_s1_readdata                     : std_logic_vector(31 downto 0); -- UART_TX_32_PO:readdata -> mm_interconnect_0:UART_TX_32_PO_s1_readdata
	signal mm_interconnect_0_uart_tx_32_po_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:UART_TX_32_PO_s1_address -> UART_TX_32_PO:address
	signal mm_interconnect_0_uart_tx_32_po_s1_write                        : std_logic;                     -- mm_interconnect_0:UART_TX_32_PO_s1_write -> mm_interconnect_0_uart_tx_32_po_s1_write:in
	signal mm_interconnect_0_uart_tx_32_po_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:UART_TX_32_PO_s1_writedata -> UART_TX_32_PO:writedata
	signal mm_interconnect_0_uart_rx_32_po_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:UART_RX_32_PO_s1_chipselect -> UART_RX_32_PO:chipselect
	signal mm_interconnect_0_uart_rx_32_po_s1_readdata                     : std_logic_vector(31 downto 0); -- UART_RX_32_PO:readdata -> mm_interconnect_0:UART_RX_32_PO_s1_readdata
	signal mm_interconnect_0_uart_rx_32_po_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:UART_RX_32_PO_s1_address -> UART_RX_32_PO:address
	signal mm_interconnect_0_uart_rx_32_po_s1_write                        : std_logic;                     -- mm_interconnect_0:UART_RX_32_PO_s1_write -> mm_interconnect_0_uart_rx_32_po_s1_write:in
	signal mm_interconnect_0_uart_rx_32_po_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:UART_RX_32_PO_s1_writedata -> UART_RX_32_PO:writedata
	signal mm_interconnect_0_uart_rx_data_reg_s1_readdata                  : std_logic_vector(31 downto 0); -- UART_RX_DATA_REG:readdata -> mm_interconnect_0:UART_RX_DATA_REG_s1_readdata
	signal mm_interconnect_0_uart_rx_data_reg_s1_address                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:UART_RX_DATA_REG_s1_address -> UART_RX_DATA_REG:address
	signal mm_interconnect_0_uart_tx_data_reg_s1_chipselect                : std_logic;                     -- mm_interconnect_0:UART_TX_DATA_REG_s1_chipselect -> UART_TX_DATA_REG:chipselect
	signal mm_interconnect_0_uart_tx_data_reg_s1_readdata                  : std_logic_vector(31 downto 0); -- UART_TX_DATA_REG:readdata -> mm_interconnect_0:UART_TX_DATA_REG_s1_readdata
	signal mm_interconnect_0_uart_tx_data_reg_s1_address                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:UART_TX_DATA_REG_s1_address -> UART_TX_DATA_REG:address
	signal mm_interconnect_0_uart_tx_data_reg_s1_write                     : std_logic;                     -- mm_interconnect_0:UART_TX_DATA_REG_s1_write -> mm_interconnect_0_uart_tx_data_reg_s1_write:in
	signal mm_interconnect_0_uart_tx_data_reg_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:UART_TX_DATA_REG_s1_writedata -> UART_TX_DATA_REG:writedata
	signal mm_interconnect_0_uart_rx_status_reg_s1_readdata                : std_logic_vector(31 downto 0); -- UART_RX_STATUS_REG:readdata -> mm_interconnect_0:UART_RX_STATUS_REG_s1_readdata
	signal mm_interconnect_0_uart_rx_status_reg_s1_address                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:UART_RX_STATUS_REG_s1_address -> UART_RX_STATUS_REG:address
	signal mm_interconnect_0_uart_tx_start_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:UART_TX_START_s1_chipselect -> UART_TX_START:chipselect
	signal mm_interconnect_0_uart_tx_start_s1_readdata                     : std_logic_vector(31 downto 0); -- UART_TX_START:readdata -> mm_interconnect_0:UART_TX_START_s1_readdata
	signal mm_interconnect_0_uart_tx_start_s1_address                      : std_logic_vector(2 downto 0);  -- mm_interconnect_0:UART_TX_START_s1_address -> UART_TX_START:address
	signal mm_interconnect_0_uart_tx_start_s1_write                        : std_logic;                     -- mm_interconnect_0:UART_TX_START_s1_write -> mm_interconnect_0_uart_tx_start_s1_write:in
	signal mm_interconnect_0_uart_tx_start_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:UART_TX_START_s1_writedata -> UART_TX_START:writedata
	signal mm_interconnect_0_control_pio_s1_readdata                       : std_logic_vector(31 downto 0); -- Control_PIO:readdata -> mm_interconnect_0:Control_PIO_s1_readdata
	signal mm_interconnect_0_control_pio_s1_address                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:Control_PIO_s1_address -> Control_PIO:address
	signal mm_interconnect_0_status_leds_pio_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:Status_LEDS_PIO_s1_chipselect -> Status_LEDS_PIO:chipselect
	signal mm_interconnect_0_status_leds_pio_s1_readdata                   : std_logic_vector(31 downto 0); -- Status_LEDS_PIO:readdata -> mm_interconnect_0:Status_LEDS_PIO_s1_readdata
	signal mm_interconnect_0_status_leds_pio_s1_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:Status_LEDS_PIO_s1_address -> Status_LEDS_PIO:address
	signal mm_interconnect_0_status_leds_pio_s1_write                      : std_logic;                     -- mm_interconnect_0:Status_LEDS_PIO_s1_write -> mm_interconnect_0_status_leds_pio_s1_write:in
	signal mm_interconnect_0_status_leds_pio_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:Status_LEDS_PIO_s1_writedata -> Status_LEDS_PIO:writedata
	signal mm_interconnect_0_dip_tx_data_pio_s1_readdata                   : std_logic_vector(31 downto 0); -- DIP_TX_Data_PIO:readdata -> mm_interconnect_0:DIP_TX_Data_PIO_s1_readdata
	signal mm_interconnect_0_dip_tx_data_pio_s1_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:DIP_TX_Data_PIO_s1_address -> DIP_TX_Data_PIO:address
	signal mm_interconnect_0_parsedloop_irq_s1_chipselect                  : std_logic;                     -- mm_interconnect_0:ParsedLoop_IRQ_s1_chipselect -> ParsedLoop_IRQ:chipselect
	signal mm_interconnect_0_parsedloop_irq_s1_readdata                    : std_logic_vector(31 downto 0); -- ParsedLoop_IRQ:readdata -> mm_interconnect_0:ParsedLoop_IRQ_s1_readdata
	signal mm_interconnect_0_parsedloop_irq_s1_address                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ParsedLoop_IRQ_s1_address -> ParsedLoop_IRQ:address
	signal mm_interconnect_0_parsedloop_irq_s1_write                       : std_logic;                     -- mm_interconnect_0:ParsedLoop_IRQ_s1_write -> mm_interconnect_0_parsedloop_irq_s1_write:in
	signal mm_interconnect_0_parsedloop_irq_s1_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:ParsedLoop_IRQ_s1_writedata -> ParsedLoop_IRQ:writedata
	signal mm_interconnect_0_uart_rx_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:UART_RX_s1_chipselect -> UART_RX:chipselect
	signal mm_interconnect_0_uart_rx_s1_readdata                           : std_logic_vector(31 downto 0); -- UART_RX:readdata -> mm_interconnect_0:UART_RX_s1_readdata
	signal mm_interconnect_0_uart_rx_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:UART_RX_s1_address -> UART_RX:address
	signal mm_interconnect_0_uart_rx_s1_write                              : std_logic;                     -- mm_interconnect_0:UART_RX_s1_write -> mm_interconnect_0_uart_rx_s1_write:in
	signal mm_interconnect_0_uart_rx_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:UART_RX_s1_writedata -> UART_RX:writedata
	signal mm_interconnect_0_uart_tx_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:UART_TX_s1_chipselect -> UART_TX:chipselect
	signal mm_interconnect_0_uart_tx_s1_readdata                           : std_logic_vector(31 downto 0); -- UART_TX:readdata -> mm_interconnect_0:UART_TX_s1_readdata
	signal mm_interconnect_0_uart_tx_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:UART_TX_s1_address -> UART_TX:address
	signal mm_interconnect_0_uart_tx_s1_write                              : std_logic;                     -- mm_interconnect_0:UART_TX_s1_write -> mm_interconnect_0_uart_tx_s1_write:in
	signal mm_interconnect_0_uart_tx_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:UART_TX_s1_writedata -> UART_TX:writedata
	signal mm_interconnect_0_start_timer_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:Start_Timer_s1_chipselect -> Start_Timer:chipselect
	signal mm_interconnect_0_start_timer_s1_readdata                       : std_logic_vector(31 downto 0); -- Start_Timer:readdata -> mm_interconnect_0:Start_Timer_s1_readdata
	signal mm_interconnect_0_start_timer_s1_address                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:Start_Timer_s1_address -> Start_Timer:address
	signal mm_interconnect_0_start_timer_s1_write                          : std_logic;                     -- mm_interconnect_0:Start_Timer_s1_write -> mm_interconnect_0_start_timer_s1_write:in
	signal mm_interconnect_0_start_timer_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:Start_Timer_s1_writedata -> Start_Timer:writedata
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- ParsedLoop_IRQ:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- UART_RX:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- UART_TX:irq -> irq_mapper:receiver3_irq
	signal nios2_gen2_0_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal nios2_gen2_0_debug_reset_request_reset                          : std_logic;                     -- nios2_gen2_0:debug_reset_request -> rst_controller:reset_in1
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_uart_tx_32_po_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_uart_tx_32_po_s1_write:inv -> UART_TX_32_PO:write_n
	signal mm_interconnect_0_uart_rx_32_po_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_uart_rx_32_po_s1_write:inv -> UART_RX_32_PO:write_n
	signal mm_interconnect_0_uart_tx_data_reg_s1_write_ports_inv           : std_logic;                     -- mm_interconnect_0_uart_tx_data_reg_s1_write:inv -> UART_TX_DATA_REG:write_n
	signal mm_interconnect_0_uart_tx_start_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_uart_tx_start_s1_write:inv -> UART_TX_START:write_n
	signal mm_interconnect_0_status_leds_pio_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_status_leds_pio_s1_write:inv -> Status_LEDS_PIO:write_n
	signal mm_interconnect_0_parsedloop_irq_s1_write_ports_inv             : std_logic;                     -- mm_interconnect_0_parsedloop_irq_s1_write:inv -> ParsedLoop_IRQ:write_n
	signal mm_interconnect_0_uart_rx_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_uart_rx_s1_write:inv -> UART_RX:write_n
	signal mm_interconnect_0_uart_tx_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_uart_tx_s1_write:inv -> UART_TX:write_n
	signal mm_interconnect_0_start_timer_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_start_timer_s1_write:inv -> Start_Timer:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Control_PIO:reset_n, DIP_TX_Data_PIO:reset_n, ParsedLoop_IRQ:reset_n, Start_Timer:reset_n, Status_LEDS_PIO:reset_n, UART_RX:reset_n, UART_RX_32_PO:reset_n, UART_RX_DATA_REG:reset_n, UART_RX_STATUS_REG:reset_n, UART_TX:reset_n, UART_TX_32_PO:reset_n, UART_TX_DATA_REG:reset_n, UART_TX_START:reset_n, nios2_gen2_0:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> jtag_uart_0:rst_n

begin

	control_pio : component NIOS2_Control_PIO
		port map (
			clk      => clk_clk,                                   --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address  => mm_interconnect_0_control_pio_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_control_pio_s1_readdata, --                    .readdata
			in_port  => control_pio_external_connection_export     -- external_connection.export
		);

	dip_tx_data_pio : component NIOS2_DIP_TX_Data_PIO
		port map (
			clk      => clk_clk,                                       --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address  => mm_interconnect_0_dip_tx_data_pio_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_dip_tx_data_pio_s1_readdata, --                    .readdata
			in_port  => dip_tx_data_pio_external_connection_export     -- external_connection.export
		);

	parsedloop_irq : component NIOS2_ParsedLoop_IRQ
		port map (
			clk        => clk_clk,                                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address    => mm_interconnect_0_parsedloop_irq_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_parsedloop_irq_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_parsedloop_irq_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_parsedloop_irq_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_parsedloop_irq_s1_readdata,        --                    .readdata
			in_port    => parsedloop_irq_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver1_irq                             --                 irq.irq
		);

	start_timer : component NIOS2_Start_Timer
		port map (
			clk        => clk_clk,                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_start_timer_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_start_timer_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_start_timer_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_start_timer_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_start_timer_s1_readdata,        --                    .readdata
			out_port   => start_timer_external_connection_export            -- external_connection.export
		);

	status_leds_pio : component NIOS2_Status_LEDS_PIO
		port map (
			clk        => clk_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => mm_interconnect_0_status_leds_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_status_leds_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_status_leds_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_status_leds_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_status_leds_pio_s1_readdata,        --                    .readdata
			out_port   => status_leds_pio_external_connection_export            -- external_connection.export
		);

	uart_rx : component NIOS2_UART_RX
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_uart_rx_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_uart_rx_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_uart_rx_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_uart_rx_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_uart_rx_s1_readdata,        --                    .readdata
			in_port    => uart_rx_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver2_irq                      --                 irq.irq
		);

	uart_rx_32_po : component NIOS2_UART_RX_32_PO
		port map (
			clk        => clk_clk,                                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => mm_interconnect_0_uart_rx_32_po_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_uart_rx_32_po_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_uart_rx_32_po_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_uart_rx_32_po_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_uart_rx_32_po_s1_readdata,        --                    .readdata
			out_port   => uart_rx_pi_external_connection_export               -- external_connection.export
		);

	uart_rx_data_reg : component NIOS2_DIP_TX_Data_PIO
		port map (
			clk      => clk_clk,                                        --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address  => mm_interconnect_0_uart_rx_data_reg_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_uart_rx_data_reg_s1_readdata, --                    .readdata
			in_port  => uart_rx_data_reg_external_connection_export     -- external_connection.export
		);

	uart_rx_status_reg : component NIOS2_UART_RX_STATUS_REG
		port map (
			clk      => clk_clk,                                          --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address  => mm_interconnect_0_uart_rx_status_reg_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_uart_rx_status_reg_s1_readdata, --                    .readdata
			in_port  => uart_rx_status_reg_external_connection_export     -- external_connection.export
		);

	uart_tx : component NIOS2_UART_RX
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_uart_tx_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_uart_tx_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_uart_tx_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_uart_tx_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_uart_tx_s1_readdata,        --                    .readdata
			in_port    => uart_tx_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver3_irq                      --                 irq.irq
		);

	uart_tx_32_po : component NIOS2_UART_RX_32_PO
		port map (
			clk        => clk_clk,                                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => mm_interconnect_0_uart_tx_32_po_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_uart_tx_32_po_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_uart_tx_32_po_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_uart_tx_32_po_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_uart_tx_32_po_s1_readdata,        --                    .readdata
			out_port   => uart_tx_po_external_connection_export               -- external_connection.export
		);

	uart_tx_data_reg : component NIOS2_UART_TX_DATA_REG
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_uart_tx_data_reg_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_uart_tx_data_reg_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_uart_tx_data_reg_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_uart_tx_data_reg_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_uart_tx_data_reg_s1_readdata,        --                    .readdata
			out_port   => uart_tx_data_reg_external_connection_export            -- external_connection.export
		);

	uart_tx_start : component NIOS2_Start_Timer
		port map (
			clk        => clk_clk,                                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => mm_interconnect_0_uart_tx_start_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_uart_tx_start_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_uart_tx_start_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_uart_tx_start_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_uart_tx_start_s1_readdata,        --                    .readdata
			out_port   => uart_tx_start_external_connection_export            -- external_connection.export
		);

	jtag_uart_0 : component NIOS2_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	nios2_gen2_0 : component NIOS2_nios2_gen2_0
		port map (
			clk                                 => clk_clk,                                                    --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_gen2_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_gen2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component NIOS2_onchip_memory2_0
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	mm_interconnect_0 : component NIOS2_mm_interconnect_0
		port map (
			clk_0_clk_clk                                  => clk_clk,                                                     --                                clk_0_clk.clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset  => rst_controller_001_reset_out_reset,                          --  jtag_uart_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                              -- nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address               => nios2_gen2_0_data_master_address,                            --                 nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest           => nios2_gen2_0_data_master_waitrequest,                        --                                         .waitrequest
			nios2_gen2_0_data_master_byteenable            => nios2_gen2_0_data_master_byteenable,                         --                                         .byteenable
			nios2_gen2_0_data_master_read                  => nios2_gen2_0_data_master_read,                               --                                         .read
			nios2_gen2_0_data_master_readdata              => nios2_gen2_0_data_master_readdata,                           --                                         .readdata
			nios2_gen2_0_data_master_readdatavalid         => nios2_gen2_0_data_master_readdatavalid,                      --                                         .readdatavalid
			nios2_gen2_0_data_master_write                 => nios2_gen2_0_data_master_write,                              --                                         .write
			nios2_gen2_0_data_master_writedata             => nios2_gen2_0_data_master_writedata,                          --                                         .writedata
			nios2_gen2_0_data_master_debugaccess           => nios2_gen2_0_data_master_debugaccess,                        --                                         .debugaccess
			nios2_gen2_0_instruction_master_address        => nios2_gen2_0_instruction_master_address,                     --          nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest    => nios2_gen2_0_instruction_master_waitrequest,                 --                                         .waitrequest
			nios2_gen2_0_instruction_master_read           => nios2_gen2_0_instruction_master_read,                        --                                         .read
			nios2_gen2_0_instruction_master_readdata       => nios2_gen2_0_instruction_master_readdata,                    --                                         .readdata
			nios2_gen2_0_instruction_master_readdatavalid  => nios2_gen2_0_instruction_master_readdatavalid,               --                                         .readdatavalid
			Control_PIO_s1_address                         => mm_interconnect_0_control_pio_s1_address,                    --                           Control_PIO_s1.address
			Control_PIO_s1_readdata                        => mm_interconnect_0_control_pio_s1_readdata,                   --                                         .readdata
			DIP_TX_Data_PIO_s1_address                     => mm_interconnect_0_dip_tx_data_pio_s1_address,                --                       DIP_TX_Data_PIO_s1.address
			DIP_TX_Data_PIO_s1_readdata                    => mm_interconnect_0_dip_tx_data_pio_s1_readdata,               --                                         .readdata
			jtag_uart_0_avalon_jtag_slave_address          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --            jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                         .write
			jtag_uart_0_avalon_jtag_slave_read             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                         .read
			jtag_uart_0_avalon_jtag_slave_readdata         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                         .readdata
			jtag_uart_0_avalon_jtag_slave_writedata        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                         .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                         .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                         .chipselect
			nios2_gen2_0_debug_mem_slave_address           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,      --             nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,        --                                         .write
			nios2_gen2_0_debug_mem_slave_read              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,         --                                         .read
			nios2_gen2_0_debug_mem_slave_readdata          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,     --                                         .readdata
			nios2_gen2_0_debug_mem_slave_writedata         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,    --                                         .writedata
			nios2_gen2_0_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,   --                                         .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,  --                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,  --                                         .debugaccess
			onchip_memory2_0_s1_address                    => mm_interconnect_0_onchip_memory2_0_s1_address,               --                      onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                      => mm_interconnect_0_onchip_memory2_0_s1_write,                 --                                         .write
			onchip_memory2_0_s1_readdata                   => mm_interconnect_0_onchip_memory2_0_s1_readdata,              --                                         .readdata
			onchip_memory2_0_s1_writedata                  => mm_interconnect_0_onchip_memory2_0_s1_writedata,             --                                         .writedata
			onchip_memory2_0_s1_byteenable                 => mm_interconnect_0_onchip_memory2_0_s1_byteenable,            --                                         .byteenable
			onchip_memory2_0_s1_chipselect                 => mm_interconnect_0_onchip_memory2_0_s1_chipselect,            --                                         .chipselect
			onchip_memory2_0_s1_clken                      => mm_interconnect_0_onchip_memory2_0_s1_clken,                 --                                         .clken
			ParsedLoop_IRQ_s1_address                      => mm_interconnect_0_parsedloop_irq_s1_address,                 --                        ParsedLoop_IRQ_s1.address
			ParsedLoop_IRQ_s1_write                        => mm_interconnect_0_parsedloop_irq_s1_write,                   --                                         .write
			ParsedLoop_IRQ_s1_readdata                     => mm_interconnect_0_parsedloop_irq_s1_readdata,                --                                         .readdata
			ParsedLoop_IRQ_s1_writedata                    => mm_interconnect_0_parsedloop_irq_s1_writedata,               --                                         .writedata
			ParsedLoop_IRQ_s1_chipselect                   => mm_interconnect_0_parsedloop_irq_s1_chipselect,              --                                         .chipselect
			Start_Timer_s1_address                         => mm_interconnect_0_start_timer_s1_address,                    --                           Start_Timer_s1.address
			Start_Timer_s1_write                           => mm_interconnect_0_start_timer_s1_write,                      --                                         .write
			Start_Timer_s1_readdata                        => mm_interconnect_0_start_timer_s1_readdata,                   --                                         .readdata
			Start_Timer_s1_writedata                       => mm_interconnect_0_start_timer_s1_writedata,                  --                                         .writedata
			Start_Timer_s1_chipselect                      => mm_interconnect_0_start_timer_s1_chipselect,                 --                                         .chipselect
			Status_LEDS_PIO_s1_address                     => mm_interconnect_0_status_leds_pio_s1_address,                --                       Status_LEDS_PIO_s1.address
			Status_LEDS_PIO_s1_write                       => mm_interconnect_0_status_leds_pio_s1_write,                  --                                         .write
			Status_LEDS_PIO_s1_readdata                    => mm_interconnect_0_status_leds_pio_s1_readdata,               --                                         .readdata
			Status_LEDS_PIO_s1_writedata                   => mm_interconnect_0_status_leds_pio_s1_writedata,              --                                         .writedata
			Status_LEDS_PIO_s1_chipselect                  => mm_interconnect_0_status_leds_pio_s1_chipselect,             --                                         .chipselect
			UART_RX_s1_address                             => mm_interconnect_0_uart_rx_s1_address,                        --                               UART_RX_s1.address
			UART_RX_s1_write                               => mm_interconnect_0_uart_rx_s1_write,                          --                                         .write
			UART_RX_s1_readdata                            => mm_interconnect_0_uart_rx_s1_readdata,                       --                                         .readdata
			UART_RX_s1_writedata                           => mm_interconnect_0_uart_rx_s1_writedata,                      --                                         .writedata
			UART_RX_s1_chipselect                          => mm_interconnect_0_uart_rx_s1_chipselect,                     --                                         .chipselect
			UART_RX_32_PO_s1_address                       => mm_interconnect_0_uart_rx_32_po_s1_address,                  --                         UART_RX_32_PO_s1.address
			UART_RX_32_PO_s1_write                         => mm_interconnect_0_uart_rx_32_po_s1_write,                    --                                         .write
			UART_RX_32_PO_s1_readdata                      => mm_interconnect_0_uart_rx_32_po_s1_readdata,                 --                                         .readdata
			UART_RX_32_PO_s1_writedata                     => mm_interconnect_0_uart_rx_32_po_s1_writedata,                --                                         .writedata
			UART_RX_32_PO_s1_chipselect                    => mm_interconnect_0_uart_rx_32_po_s1_chipselect,               --                                         .chipselect
			UART_RX_DATA_REG_s1_address                    => mm_interconnect_0_uart_rx_data_reg_s1_address,               --                      UART_RX_DATA_REG_s1.address
			UART_RX_DATA_REG_s1_readdata                   => mm_interconnect_0_uart_rx_data_reg_s1_readdata,              --                                         .readdata
			UART_RX_STATUS_REG_s1_address                  => mm_interconnect_0_uart_rx_status_reg_s1_address,             --                    UART_RX_STATUS_REG_s1.address
			UART_RX_STATUS_REG_s1_readdata                 => mm_interconnect_0_uart_rx_status_reg_s1_readdata,            --                                         .readdata
			UART_TX_s1_address                             => mm_interconnect_0_uart_tx_s1_address,                        --                               UART_TX_s1.address
			UART_TX_s1_write                               => mm_interconnect_0_uart_tx_s1_write,                          --                                         .write
			UART_TX_s1_readdata                            => mm_interconnect_0_uart_tx_s1_readdata,                       --                                         .readdata
			UART_TX_s1_writedata                           => mm_interconnect_0_uart_tx_s1_writedata,                      --                                         .writedata
			UART_TX_s1_chipselect                          => mm_interconnect_0_uart_tx_s1_chipselect,                     --                                         .chipselect
			UART_TX_32_PO_s1_address                       => mm_interconnect_0_uart_tx_32_po_s1_address,                  --                         UART_TX_32_PO_s1.address
			UART_TX_32_PO_s1_write                         => mm_interconnect_0_uart_tx_32_po_s1_write,                    --                                         .write
			UART_TX_32_PO_s1_readdata                      => mm_interconnect_0_uart_tx_32_po_s1_readdata,                 --                                         .readdata
			UART_TX_32_PO_s1_writedata                     => mm_interconnect_0_uart_tx_32_po_s1_writedata,                --                                         .writedata
			UART_TX_32_PO_s1_chipselect                    => mm_interconnect_0_uart_tx_32_po_s1_chipselect,               --                                         .chipselect
			UART_TX_DATA_REG_s1_address                    => mm_interconnect_0_uart_tx_data_reg_s1_address,               --                      UART_TX_DATA_REG_s1.address
			UART_TX_DATA_REG_s1_write                      => mm_interconnect_0_uart_tx_data_reg_s1_write,                 --                                         .write
			UART_TX_DATA_REG_s1_readdata                   => mm_interconnect_0_uart_tx_data_reg_s1_readdata,              --                                         .readdata
			UART_TX_DATA_REG_s1_writedata                  => mm_interconnect_0_uart_tx_data_reg_s1_writedata,             --                                         .writedata
			UART_TX_DATA_REG_s1_chipselect                 => mm_interconnect_0_uart_tx_data_reg_s1_chipselect,            --                                         .chipselect
			UART_TX_START_s1_address                       => mm_interconnect_0_uart_tx_start_s1_address,                  --                         UART_TX_START_s1.address
			UART_TX_START_s1_write                         => mm_interconnect_0_uart_tx_start_s1_write,                    --                                         .write
			UART_TX_START_s1_readdata                      => mm_interconnect_0_uart_tx_start_s1_readdata,                 --                                         .readdata
			UART_TX_START_s1_writedata                     => mm_interconnect_0_uart_tx_start_s1_writedata,                --                                         .writedata
			UART_TX_START_s1_chipselect                    => mm_interconnect_0_uart_tx_start_s1_chipselect                --                                         .chipselect
		);

	irq_mapper : component NIOS2_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component nios2_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_001 : component nios2_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_uart_tx_32_po_s1_write_ports_inv <= not mm_interconnect_0_uart_tx_32_po_s1_write;

	mm_interconnect_0_uart_rx_32_po_s1_write_ports_inv <= not mm_interconnect_0_uart_rx_32_po_s1_write;

	mm_interconnect_0_uart_tx_data_reg_s1_write_ports_inv <= not mm_interconnect_0_uart_tx_data_reg_s1_write;

	mm_interconnect_0_uart_tx_start_s1_write_ports_inv <= not mm_interconnect_0_uart_tx_start_s1_write;

	mm_interconnect_0_status_leds_pio_s1_write_ports_inv <= not mm_interconnect_0_status_leds_pio_s1_write;

	mm_interconnect_0_parsedloop_irq_s1_write_ports_inv <= not mm_interconnect_0_parsedloop_irq_s1_write;

	mm_interconnect_0_uart_rx_s1_write_ports_inv <= not mm_interconnect_0_uart_rx_s1_write;

	mm_interconnect_0_uart_tx_s1_write_ports_inv <= not mm_interconnect_0_uart_tx_s1_write;

	mm_interconnect_0_start_timer_s1_write_ports_inv <= not mm_interconnect_0_start_timer_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of NIOS2
